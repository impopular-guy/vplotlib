module vplotlib

pub const (
	version = '0.1.1'
)
