module vplotlib

pub fn version() string {
	return "0.0.0"
}
